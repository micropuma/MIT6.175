function
    
endfunction